typedef enum {
  NONE = 0,
  LEFT, RIGHT, DOWN, DROP,
  HOLD, ROTATE, ROTATE_REV, BAR
} control_type;
